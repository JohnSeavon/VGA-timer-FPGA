LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DE0_NANO IS
    PORT ( 
		CLOCK_50 : IN STD_LOGIC;
		Reset		: IN STD_LOGIC;
		VGA_HS	: OUT STD_LOGIC;		
		VGA_VS	: OUT STD_LOGIC;
		VGA_R		: OUT STD_LOGIC_VECTOR (0 TO 3);
		VGA_G		: OUT STD_LOGIC_VECTOR (0 TO 3);
		VGA_B		: OUT STD_LOGIC_VECTOR (0 TO 3));
END DE0_NANO;

ARCHITECTURE arch OF DE0_NANO IS

COMPONENT vga_clock IS
	PORT(
		RESET : IN STD_LOGIC;
		F_CLOCK : IN STD_LOGIC;
		F_HSYNC : OUT STD_LOGIC;
		F_VSYNC : OUT STD_LOGIC;
		F_ROW : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		F_COLUMN : OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
		F_DISP_ENABLE : OUT STD_LOGIC
	);
END COMPONENT vga_clock;

COMPONENT PixelGen IS
	PORT(
		RESET : IN STD_LOGIC;
		F_CLOCK : IN STD_LOGIC;
		F_ON : IN STD_LOGIC;
		F_ROW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		F_COLUMN : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		R_OUT : OUT STD_LOGIC_VECTOR (0 TO 3); -- Componente R
		G_OUT : OUT STD_LOGIC_VECTOR (0 To 3); -- Componente G
		B_OUT : OUT STD_LOGIC_VECTOR (0 TO 3)-- Componente B
	);
END COMPONENT PixelGen;

--Índice da linha/coluna atual
SIGNAL CURRENT_ROW : STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL CURRENT_COLUMN : STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL DISP_ENABLE : STD_LOGIC;

SIGNAL HSYNC: STD_LOGIC;
SIGNAL VSYNC: STD_LOGIC;
SIGNAL Rp: STD_LOGIC_VECTOR (0 to 3);
SIGNAL Gp: STD_LOGIC_VECTOR (0 to 3);
SIGNAL Bp: STD_LOGIC_VECTOR (0 to 3);

BEGIN

	--Módulo de sincronismo
	VGA : vga_clock PORT MAP(
				RESET => RESET,
				F_CLOCK => CLOCK_50, 
				F_HSYNC => VGA_HS, 
				F_VSYNC => VGA_VS, 
				F_ROW => CURRENT_ROW,
				F_COLUMN => CURRENT_COLUMN,
				F_DISP_ENABLE => DISP_ENABLE);

	--Módulo para gerar os pixels
	PIXELS : PixelGen PORT MAP(
				RESET => RESET,
				F_CLOCK => CLOCK_50, 
				F_ON => DISP_ENABLE,
				F_ROW => CURRENT_ROW,
				F_COLUMN => CURRENT_COLUMN,
				R_OUT => Rp,
				G_OUT => Gp,
				B_OUT => Bp);
	
	PROCESS(CLOCK_50)
 BEGIN
         IF CLOCK_50'EVENT AND CLOCK_50='1' THEN
 
 VGA_VS <= VSYNC;
 VGA_HS <= HSYNC;
 VGA_R <= Rp; 
 VGA_G <= Gp;
 VGA_B <= Bp;
 
 END IF;
 END PROCESS;
END arch;